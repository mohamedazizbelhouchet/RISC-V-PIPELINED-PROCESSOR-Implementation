module instruction_memory( 
	 input  clk,
    input  [31:0] PCF,
	 input  write_enable,
	 input  [31:0] data_in,
    output wire [31:0] RD );
	 
	 reg [7:0] mem [1023:0]; /*= {  {8'h00}, {8'h11}, {8'h22}, {8'h33}, {8'h44}, {8'h55}, {8'h66}, {8'h77},
              {8'h88}, {8'h99}, {8'hAA}, {8'hBB}, {8'hCC}, {8'hDD}, {8'hEE}, {8'hFF} ,
            // Repeat as needed
            { {1024-16{8'h00}} } }  ;*/
	 reg [31:0] temp_data_out;
	 always @(*) begin 
			temp_data_out = {mem[PCF+3],mem[PCF+2],mem[PCF+1],mem[PCF]};
		end
		 

    // Assign the temporary variable to the output
    assign RD = temp_data_out;
     
	 always @(posedge clk) begin
        if (write_enable) 
            mem[PCF] <= data_in[7:0];
				mem[PCF+1] <= data_in[15:8];
				mem[PCF+2] <= data_in[23:16];
				mem[PCF+3] <= data_in[31:24];		
        end

    initial begin
    mem[ 0 ]=8'd 0  ;
mem[ 1 ]=8'd 1  ;
mem[ 2 ]=8'd 2  ;
mem[ 3 ]=8'd 3  ;
mem[ 4 ]=8'd 4  ;
mem[ 5 ]=8'd 5  ;
mem[ 6 ]=8'd 6  ;
mem[ 7 ]=8'd 7  ;
mem[ 8 ]=8'd 8  ;
mem[ 9 ]=8'd 9  ;
mem[ 10 ]=8'd 10  ;
mem[ 11 ]=8'd 11  ;
mem[ 12 ]=8'd 12  ;
mem[ 13 ]=8'd 13  ;
mem[ 14 ]=8'd 14  ;
mem[ 15 ]=8'd 15  ;
mem[ 16 ]=8'd 16  ;
mem[ 17 ]=8'd 17  ;
mem[ 18 ]=8'd 18  ;
mem[ 19 ]=8'd 19  ;
mem[ 20 ]=8'd 20  ;
mem[ 21 ]=8'd 21  ;
mem[ 22 ]=8'd 22  ;
mem[ 23 ]=8'd 23  ;
mem[ 24 ]=8'd 24  ;
mem[ 25 ]=8'd 25  ;
mem[ 26 ]=8'd 26  ;
mem[ 27 ]=8'd 27  ;
mem[ 28 ]=8'd 28  ;
mem[ 29 ]=8'd 29  ;
mem[ 30 ]=8'd 30  ;
mem[ 31 ]=8'd 31  ;
mem[ 32 ]=8'd 32  ;
mem[ 33 ]=8'd 33  ;
mem[ 34 ]=8'd 34  ;
mem[ 35 ]=8'd 35  ;
mem[ 36 ]=8'd 36  ;
mem[ 37 ]=8'd 37  ;
mem[ 38 ]=8'd 38  ;
mem[ 39 ]=8'd 39  ;
mem[ 40 ]=8'd 40  ;
mem[ 41 ]=8'd 41  ;
mem[ 42 ]=8'd 42  ;
mem[ 43 ]=8'd 43  ;
mem[ 44 ]=8'd 44  ;
mem[ 45 ]=8'd 45  ;
mem[ 46 ]=8'd 46  ;
mem[ 47 ]=8'd 47  ;
mem[ 48 ]=8'd 48  ;
mem[ 49 ]=8'd 49  ;
mem[ 50 ]=8'd 50  ;
mem[ 51 ]=8'd 51  ;
mem[ 52 ]=8'd 52  ;
mem[ 53 ]=8'd 53  ;
mem[ 54 ]=8'd 54  ;
mem[ 55 ]=8'd 55  ;
mem[ 56 ]=8'd 56  ;
mem[ 57 ]=8'd 57  ;
mem[ 58 ]=8'd 58  ;
mem[ 59 ]=8'd 59  ;
mem[ 60 ]=8'd 60  ;
mem[ 61 ]=8'd 61  ;
mem[ 62 ]=8'd 62  ;
mem[ 63 ]=8'd 63  ;
mem[ 64 ]=8'd 64  ;
mem[ 65 ]=8'd 65  ;
mem[ 66 ]=8'd 66  ;
mem[ 67 ]=8'd 67  ;
mem[ 68 ]=8'd 68  ;
mem[ 69 ]=8'd 69  ;
mem[ 70 ]=8'd 70  ;
mem[ 71 ]=8'd 71  ;
mem[ 72 ]=8'd 72  ;
mem[ 73 ]=8'd 73  ;
mem[ 74 ]=8'd 74  ;
mem[ 75 ]=8'd 75  ;
mem[ 76 ]=8'd 76  ;
mem[ 77 ]=8'd 77  ;
mem[ 78 ]=8'd 78  ;
mem[ 79 ]=8'd 79  ;
mem[ 80 ]=8'd 80  ;
mem[ 81 ]=8'd 81  ;
mem[ 82 ]=8'd 82  ;
mem[ 83 ]=8'd 83  ;
mem[ 84 ]=8'd 84  ;
mem[ 85 ]=8'd 85  ;
mem[ 86 ]=8'd 86  ;
mem[ 87 ]=8'd 87  ;
mem[ 88 ]=8'd 88  ;
mem[ 89 ]=8'd 89  ;
mem[ 90 ]=8'd 90  ;
mem[ 91 ]=8'd 91  ;
mem[ 92 ]=8'd 92  ;
mem[ 93 ]=8'd 93  ;
mem[ 94 ]=8'd 94  ;
mem[ 95 ]=8'd 95  ;
mem[ 96 ]=8'd 96  ;
mem[ 97 ]=8'd 97  ;
mem[ 98 ]=8'd 98  ;
mem[ 99 ]=8'd 99  ;
mem[ 100 ]=8'd 100  ;
mem[ 101 ]=8'd 101  ;
mem[ 102 ]=8'd 102  ;
mem[ 103 ]=8'd 103  ;
mem[ 104 ]=8'd 104  ;
mem[ 105 ]=8'd 105  ;
mem[ 106 ]=8'd 106  ;
mem[ 107 ]=8'd 107  ;
mem[ 108 ]=8'd 108  ;
mem[ 109 ]=8'd 109  ;
mem[ 110 ]=8'd 110  ;
mem[ 111 ]=8'd 111  ;
mem[ 112 ]=8'd 112  ;
mem[ 113 ]=8'd 113  ;
mem[ 114 ]=8'd 114  ;
mem[ 115 ]=8'd 115  ;
mem[ 116 ]=8'd 116  ;
mem[ 117 ]=8'd 117  ;
mem[ 118 ]=8'd 118  ;
mem[ 119 ]=8'd 119  ;
mem[ 120 ]=8'd 120  ;
mem[ 121 ]=8'd 121  ;
mem[ 122 ]=8'd 122  ;
mem[ 123 ]=8'd 123  ;
mem[ 124 ]=8'd 124  ;
mem[ 125 ]=8'd 125  ;
mem[ 126 ]=8'd 126  ;
mem[ 127 ]=8'd 127  ;
mem[ 128 ]=8'd 128  ;
mem[ 129 ]=8'd 129  ;
mem[ 130 ]=8'd 130  ;
mem[ 131 ]=8'd 131  ;
mem[ 132 ]=8'd 132  ;
mem[ 133 ]=8'd 133  ;
mem[ 134 ]=8'd 134  ;
mem[ 135 ]=8'd 135  ;
mem[ 136 ]=8'd 136  ;
mem[ 137 ]=8'd 137  ;
mem[ 138 ]=8'd 138  ;
mem[ 139 ]=8'd 139  ;
mem[ 140 ]=8'd 140  ;
mem[ 141 ]=8'd 141  ;
mem[ 142 ]=8'd 142  ;
mem[ 143 ]=8'd 143  ;
mem[ 144 ]=8'd 144  ;
mem[ 145 ]=8'd 145  ;
mem[ 146 ]=8'd 146  ;
mem[ 147 ]=8'd 147  ;
mem[ 148 ]=8'd 148  ;
mem[ 149 ]=8'd 149  ;
mem[ 150 ]=8'd 150  ;
mem[ 151 ]=8'd 151  ;
mem[ 152 ]=8'd 152  ;
mem[ 153 ]=8'd 153  ;
mem[ 154 ]=8'd 154  ;
mem[ 155 ]=8'd 155  ;
mem[ 156 ]=8'd 156  ;
mem[ 157 ]=8'd 157  ;
mem[ 158 ]=8'd 158  ;
mem[ 159 ]=8'd 159  ;
mem[ 160 ]=8'd 160  ;
mem[ 161 ]=8'd 161  ;
mem[ 162 ]=8'd 162  ;
mem[ 163 ]=8'd 163  ;
mem[ 164 ]=8'd 164  ;
mem[ 165 ]=8'd 165  ;
mem[ 166 ]=8'd 166  ;
mem[ 167 ]=8'd 167  ;
mem[ 168 ]=8'd 168  ;
mem[ 169 ]=8'd 169  ;
mem[ 170 ]=8'd 170  ;
mem[ 171 ]=8'd 171  ;
mem[ 172 ]=8'd 172  ;
mem[ 173 ]=8'd 173  ;
mem[ 174 ]=8'd 174  ;
mem[ 175 ]=8'd 175  ;
mem[ 176 ]=8'd 176  ;
mem[ 177 ]=8'd 177  ;
mem[ 178 ]=8'd 178  ;
mem[ 179 ]=8'd 179  ;
mem[ 180 ]=8'd 180  ;
mem[ 181 ]=8'd 181  ;
mem[ 182 ]=8'd 182  ;
mem[ 183 ]=8'd 183  ;
mem[ 184 ]=8'd 184  ;
mem[ 185 ]=8'd 185  ;
mem[ 186 ]=8'd 186  ;
mem[ 187 ]=8'd 187  ;
mem[ 188 ]=8'd 188  ;
mem[ 189 ]=8'd 189  ;
mem[ 190 ]=8'd 190  ;
mem[ 191 ]=8'd 191  ;
mem[ 192 ]=8'd 192  ;
mem[ 193 ]=8'd 193  ;
mem[ 194 ]=8'd 194  ;
mem[ 195 ]=8'd 195  ;
mem[ 196 ]=8'd 196  ;
mem[ 197 ]=8'd 197  ;
mem[ 198 ]=8'd 198  ;
mem[ 199 ]=8'd 199  ;
mem[ 200 ]=8'd 200  ;
mem[ 201 ]=8'd 201  ;
mem[ 202 ]=8'd 202  ;
mem[ 203 ]=8'd 203  ;
mem[ 204 ]=8'd 204  ;
mem[ 205 ]=8'd 205  ;
mem[ 206 ]=8'd 206  ;
mem[ 207 ]=8'd 207  ;
mem[ 208 ]=8'd 208  ;
mem[ 209 ]=8'd 209  ;
mem[ 210 ]=8'd 210  ;
mem[ 211 ]=8'd 211  ;
mem[ 212 ]=8'd 212  ;
mem[ 213 ]=8'd 213  ;
mem[ 214 ]=8'd 214  ;
mem[ 215 ]=8'd 215  ;
mem[ 216 ]=8'd 216  ;
mem[ 217 ]=8'd 217  ;
mem[ 218 ]=8'd 218  ;
mem[ 219 ]=8'd 219  ;
mem[ 220 ]=8'd 220  ;
mem[ 221 ]=8'd 221  ;
mem[ 222 ]=8'd 222  ;
mem[ 223 ]=8'd 223  ;
mem[ 224 ]=8'd 224  ;
mem[ 225 ]=8'd 225  ;
mem[ 226 ]=8'd 226  ;
mem[ 227 ]=8'd 227  ;
mem[ 228 ]=8'd 228  ;
mem[ 229 ]=8'd 229  ;
mem[ 230 ]=8'd 230  ;
mem[ 231 ]=8'd 231  ;
mem[ 232 ]=8'd 232  ;
mem[ 233 ]=8'd 233  ;
mem[ 234 ]=8'd 234  ;
mem[ 235 ]=8'd 235  ;
mem[ 236 ]=8'd 236  ;
mem[ 237 ]=8'd 237  ;
mem[ 238 ]=8'd 238  ;
mem[ 239 ]=8'd 239  ;
mem[ 240 ]=8'd 240  ;
mem[ 241 ]=8'd 241  ;
mem[ 242 ]=8'd 242  ;
mem[ 243 ]=8'd 243  ;
mem[ 244 ]=8'd 244  ;
mem[ 245 ]=8'd 245  ;
mem[ 246 ]=8'd 246  ;
mem[ 247 ]=8'd 247  ;
mem[ 248 ]=8'd 248  ;
mem[ 249 ]=8'd 249  ;
mem[ 250 ]=8'd 250  ;
mem[ 251 ]=8'd 251  ;
mem[ 252 ]=8'd 252  ;
mem[ 253 ]=8'd 253  ;
mem[ 254 ]=8'd 254  ;
mem[ 255 ]=8'd 255  ;
mem[ 256 ]=8'd 256  ;
mem[ 257 ]=8'd 257  ;
mem[ 258 ]=8'd 258  ;
mem[ 259 ]=8'd 259  ;
mem[ 260 ]=8'd 260  ;
mem[ 261 ]=8'd 261  ;
mem[ 262 ]=8'd 262  ;
mem[ 263 ]=8'd 263  ;
mem[ 264 ]=8'd 264  ;
mem[ 265 ]=8'd 265  ;
mem[ 266 ]=8'd 266  ;
mem[ 267 ]=8'd 267  ;
mem[ 268 ]=8'd 268  ;
mem[ 269 ]=8'd 269  ;
mem[ 270 ]=8'd 270  ;
mem[ 271 ]=8'd 271  ;
mem[ 272 ]=8'd 272  ;
mem[ 273 ]=8'd 273  ;
mem[ 274 ]=8'd 274  ;
mem[ 275 ]=8'd 275  ;
mem[ 276 ]=8'd 276  ;
mem[ 277 ]=8'd 277  ;
mem[ 278 ]=8'd 278  ;
mem[ 279 ]=8'd 279  ;
mem[ 280 ]=8'd 280  ;
mem[ 281 ]=8'd 281  ;
mem[ 282 ]=8'd 282  ;
mem[ 283 ]=8'd 283  ;
mem[ 284 ]=8'd 284  ;
mem[ 285 ]=8'd 285  ;
mem[ 286 ]=8'd 286  ;
mem[ 287 ]=8'd 287  ;
mem[ 288 ]=8'd 288  ;
mem[ 289 ]=8'd 289  ;
mem[ 290 ]=8'd 290  ;
mem[ 291 ]=8'd 291  ;
mem[ 292 ]=8'd 292  ;
mem[ 293 ]=8'd 293  ;
mem[ 294 ]=8'd 294  ;
mem[ 295 ]=8'd 295  ;
mem[ 296 ]=8'd 296  ;
mem[ 297 ]=8'd 297  ;
mem[ 298 ]=8'd 298  ;
mem[ 299 ]=8'd 299  ;
mem[ 300 ]=8'd 300  ;
mem[ 301 ]=8'd 301  ;
mem[ 302 ]=8'd 302  ;
mem[ 303 ]=8'd 303  ;
mem[ 304 ]=8'd 304  ;
mem[ 305 ]=8'd 305  ;
mem[ 306 ]=8'd 306  ;
mem[ 307 ]=8'd 307  ;
mem[ 308 ]=8'd 308  ;
mem[ 309 ]=8'd 309  ;
mem[ 310 ]=8'd 310  ;
mem[ 311 ]=8'd 311  ;
mem[ 312 ]=8'd 312  ;
mem[ 313 ]=8'd 313  ;
mem[ 314 ]=8'd 314  ;
mem[ 315 ]=8'd 315  ;
mem[ 316 ]=8'd 316  ;
mem[ 317 ]=8'd 317  ;
mem[ 318 ]=8'd 318  ;
mem[ 319 ]=8'd 319  ;
mem[ 320 ]=8'd 320  ;
mem[ 321 ]=8'd 321  ;
mem[ 322 ]=8'd 322  ;
mem[ 323 ]=8'd 323  ;
mem[ 324 ]=8'd 324  ;
mem[ 325 ]=8'd 325  ;
mem[ 326 ]=8'd 326  ;
mem[ 327 ]=8'd 327  ;
mem[ 328 ]=8'd 328  ;
mem[ 329 ]=8'd 329  ;
mem[ 330 ]=8'd 330  ;
mem[ 331 ]=8'd 331  ;
mem[ 332 ]=8'd 332  ;
mem[ 333 ]=8'd 333  ;
mem[ 334 ]=8'd 334  ;
mem[ 335 ]=8'd 335  ;
mem[ 336 ]=8'd 336  ;
mem[ 337 ]=8'd 337  ;
mem[ 338 ]=8'd 338  ;
mem[ 339 ]=8'd 339  ;
mem[ 340 ]=8'd 340  ;
mem[ 341 ]=8'd 341  ;
mem[ 342 ]=8'd 342  ;
mem[ 343 ]=8'd 343  ;
mem[ 344 ]=8'd 344  ;
mem[ 345 ]=8'd 345  ;
mem[ 346 ]=8'd 346  ;
mem[ 347 ]=8'd 347  ;
mem[ 348 ]=8'd 348  ;
mem[ 349 ]=8'd 349  ;
mem[ 350 ]=8'd 350  ;
mem[ 351 ]=8'd 351  ;
mem[ 352 ]=8'd 352  ;
mem[ 353 ]=8'd 353  ;
mem[ 354 ]=8'd 354  ;
mem[ 355 ]=8'd 355  ;
mem[ 356 ]=8'd 356  ;
mem[ 357 ]=8'd 357  ;
mem[ 358 ]=8'd 358  ;
mem[ 359 ]=8'd 359  ;
mem[ 360 ]=8'd 360  ;
mem[ 361 ]=8'd 361  ;
mem[ 362 ]=8'd 362  ;
mem[ 363 ]=8'd 363  ;
mem[ 364 ]=8'd 364  ;
mem[ 365 ]=8'd 365  ;
mem[ 366 ]=8'd 366  ;
mem[ 367 ]=8'd 367  ;
mem[ 368 ]=8'd 368  ;
mem[ 369 ]=8'd 369  ;
mem[ 370 ]=8'd 370  ;
mem[ 371 ]=8'd 371  ;
mem[ 372 ]=8'd 372  ;
mem[ 373 ]=8'd 373  ;
mem[ 374 ]=8'd 374  ;
mem[ 375 ]=8'd 375  ;
mem[ 376 ]=8'd 376  ;
mem[ 377 ]=8'd 377  ;
mem[ 378 ]=8'd 378  ;
mem[ 379 ]=8'd 379  ;
mem[ 380 ]=8'd 380  ;
mem[ 381 ]=8'd 381  ;
mem[ 382 ]=8'd 382  ;
mem[ 383 ]=8'd 383  ;
mem[ 384 ]=8'd 384  ;
mem[ 385 ]=8'd 385  ;
mem[ 386 ]=8'd 386  ;
mem[ 387 ]=8'd 387  ;
mem[ 388 ]=8'd 388  ;
mem[ 389 ]=8'd 389  ;
mem[ 390 ]=8'd 390  ;
mem[ 391 ]=8'd 391  ;
mem[ 392 ]=8'd 392  ;
mem[ 393 ]=8'd 393  ;
mem[ 394 ]=8'd 394  ;
mem[ 395 ]=8'd 395  ;
mem[ 396 ]=8'd 396  ;
mem[ 397 ]=8'd 397  ;
mem[ 398 ]=8'd 398  ;
mem[ 399 ]=8'd 399  ;
mem[ 400 ]=8'd 400  ;
mem[ 401 ]=8'd 401  ;
mem[ 402 ]=8'd 402  ;
mem[ 403 ]=8'd 403  ;
mem[ 404 ]=8'd 404  ;
mem[ 405 ]=8'd 405  ;
mem[ 406 ]=8'd 406  ;
mem[ 407 ]=8'd 407  ;
mem[ 408 ]=8'd 408  ;
mem[ 409 ]=8'd 409  ;
mem[ 410 ]=8'd 410  ;
mem[ 411 ]=8'd 411  ;
mem[ 412 ]=8'd 412  ;
mem[ 413 ]=8'd 413  ;
mem[ 414 ]=8'd 414  ;
mem[ 415 ]=8'd 415  ;
mem[ 416 ]=8'd 416  ;
mem[ 417 ]=8'd 417  ;
mem[ 418 ]=8'd 418  ;
mem[ 419 ]=8'd 419  ;
mem[ 420 ]=8'd 420  ;
mem[ 421 ]=8'd 421  ;
mem[ 422 ]=8'd 422  ;
mem[ 423 ]=8'd 423  ;
mem[ 424 ]=8'd 424  ;
mem[ 425 ]=8'd 425  ;
mem[ 426 ]=8'd 426  ;
mem[ 427 ]=8'd 427  ;
mem[ 428 ]=8'd 428  ;
mem[ 429 ]=8'd 429  ;
mem[ 430 ]=8'd 430  ;
mem[ 431 ]=8'd 431  ;
mem[ 432 ]=8'd 432  ;
mem[ 433 ]=8'd 433  ;
mem[ 434 ]=8'd 434  ;
mem[ 435 ]=8'd 435  ;
mem[ 436 ]=8'd 436  ;
mem[ 437 ]=8'd 437  ;
mem[ 438 ]=8'd 438  ;
mem[ 439 ]=8'd 439  ;
mem[ 440 ]=8'd 440  ;
mem[ 441 ]=8'd 441  ;
mem[ 442 ]=8'd 442  ;
mem[ 443 ]=8'd 443  ;
mem[ 444 ]=8'd 444  ;
mem[ 445 ]=8'd 445  ;
mem[ 446 ]=8'd 446  ;
mem[ 447 ]=8'd 447  ;
mem[ 448 ]=8'd 448  ;
mem[ 449 ]=8'd 449  ;
mem[ 450 ]=8'd 450  ;
mem[ 451 ]=8'd 451  ;
mem[ 452 ]=8'd 452  ;
mem[ 453 ]=8'd 453  ;
mem[ 454 ]=8'd 454  ;
mem[ 455 ]=8'd 455  ;
mem[ 456 ]=8'd 456  ;
mem[ 457 ]=8'd 457  ;
mem[ 458 ]=8'd 458  ;
mem[ 459 ]=8'd 459  ;
mem[ 460 ]=8'd 460  ;
mem[ 461 ]=8'd 461  ;
mem[ 462 ]=8'd 462  ;
mem[ 463 ]=8'd 463  ;
mem[ 464 ]=8'd 464  ;
mem[ 465 ]=8'd 465  ;
mem[ 466 ]=8'd 466  ;
mem[ 467 ]=8'd 467  ;
mem[ 468 ]=8'd 468  ;
mem[ 469 ]=8'd 469  ;
mem[ 470 ]=8'd 470  ;
mem[ 471 ]=8'd 471  ;
mem[ 472 ]=8'd 472  ;
mem[ 473 ]=8'd 473  ;
mem[ 474 ]=8'd 474  ;
mem[ 475 ]=8'd 475  ;
mem[ 476 ]=8'd 476  ;
mem[ 477 ]=8'd 477  ;
mem[ 478 ]=8'd 478  ;
mem[ 479 ]=8'd 479  ;
mem[ 480 ]=8'd 480  ;
mem[ 481 ]=8'd 481  ;
mem[ 482 ]=8'd 482  ;
mem[ 483 ]=8'd 483  ;
mem[ 484 ]=8'd 484  ;
mem[ 485 ]=8'd 485  ;
mem[ 486 ]=8'd 486  ;
mem[ 487 ]=8'd 487  ;
mem[ 488 ]=8'd 488  ;
mem[ 489 ]=8'd 489  ;
mem[ 490 ]=8'd 490  ;
mem[ 491 ]=8'd 491  ;
mem[ 492 ]=8'd 492  ;
mem[ 493 ]=8'd 493  ;
mem[ 494 ]=8'd 494  ;
mem[ 495 ]=8'd 495  ;
mem[ 496 ]=8'd 496  ;
mem[ 497 ]=8'd 497  ;
mem[ 498 ]=8'd 498  ;
mem[ 499 ]=8'd 499  ;
mem[ 500 ]=8'd 500  ;
mem[ 501 ]=8'd 501  ;
mem[ 502 ]=8'd 502  ;
mem[ 503 ]=8'd 503  ;
mem[ 504 ]=8'd 504  ;
mem[ 505 ]=8'd 505  ;
mem[ 506 ]=8'd 506  ;
mem[ 507 ]=8'd 507  ;
mem[ 508 ]=8'd 508  ;
mem[ 509 ]=8'd 509  ;
mem[ 510 ]=8'd 510  ;
mem[ 511 ]=8'd 511  ;
mem[ 512 ]=8'd 512  ;
mem[ 513 ]=8'd 513  ;
mem[ 514 ]=8'd 514  ;
mem[ 515 ]=8'd 515  ;
mem[ 516 ]=8'd 516  ;
mem[ 517 ]=8'd 517  ;
mem[ 518 ]=8'd 518  ;
mem[ 519 ]=8'd 519  ;
mem[ 520 ]=8'd 520  ;
mem[ 521 ]=8'd 521  ;
mem[ 522 ]=8'd 522  ;
mem[ 523 ]=8'd 523  ;
mem[ 524 ]=8'd 524  ;
mem[ 525 ]=8'd 525  ;
mem[ 526 ]=8'd 526  ;
mem[ 527 ]=8'd 527  ;
mem[ 528 ]=8'd 528  ;
mem[ 529 ]=8'd 529  ;
mem[ 530 ]=8'd 530  ;
mem[ 531 ]=8'd 531  ;mem[ 532 ]=8'd 532  ;
mem[ 533 ]=8'd 533  ;
mem[ 534 ]=8'd 534  ;
mem[ 535 ]=8'd 535  ;
mem[ 536 ]=8'd 536  ;
mem[ 537 ]=8'd 537  ;
mem[ 538 ]=8'd 538  ;
mem[ 539 ]=8'd 539  ;
mem[ 540 ]=8'd 540  ;
mem[ 541 ]=8'd 541  ;
mem[ 542 ]=8'd 542  ;
mem[ 543 ]=8'd 543  ;
mem[ 544 ]=8'd 544  ;
mem[ 545 ]=8'd 545  ;
mem[ 546 ]=8'd 546  ;
mem[ 547 ]=8'd 547  ;
mem[ 548 ]=8'd 548  ;
mem[ 549 ]=8'd 549  ;
mem[ 550 ]=8'd 550  ;
mem[ 551 ]=8'd 551  ;
mem[ 552 ]=8'd 552  ;
mem[ 553 ]=8'd 553  ;
mem[ 554 ]=8'd 554  ;
mem[ 555 ]=8'd 555  ;
mem[ 556 ]=8'd 556  ;
mem[ 557 ]=8'd 557  ;
mem[ 558 ]=8'd 558  ;
mem[ 559 ]=8'd 559  ;
mem[ 560 ]=8'd 560  ;
mem[ 561 ]=8'd 561  ;
mem[ 562 ]=8'd 562  ;
mem[ 563 ]=8'd 563  ;
mem[ 564 ]=8'd 564  ;
mem[ 565 ]=8'd 565  ;
mem[ 566 ]=8'd 566  ;
mem[ 567 ]=8'd 567  ;
mem[ 568 ]=8'd 568  ;
mem[ 569 ]=8'd 569  ;
mem[ 570 ]=8'd 570  ;
mem[ 571 ]=8'd 571  ;
mem[ 572 ]=8'd 572  ;
mem[ 573 ]=8'd 573  ;
mem[ 574 ]=8'd 574  ;
mem[ 575 ]=8'd 575  ;
mem[ 576 ]=8'd 576  ;
mem[ 577 ]=8'd 577  ;
mem[ 578 ]=8'd 578  ;
mem[ 579 ]=8'd 579  ;
mem[ 580 ]=8'd 580  ;
mem[ 581 ]=8'd 581  ;
mem[ 582 ]=8'd 582  ;
mem[ 583 ]=8'd 583  ;
mem[ 584 ]=8'd 584  ;
mem[ 585 ]=8'd 585  ;
mem[ 586 ]=8'd 586  ;
mem[ 587 ]=8'd 587  ;
mem[ 588 ]=8'd 588  ;
mem[ 589 ]=8'd 589  ;
mem[ 590 ]=8'd 590  ;
mem[ 591 ]=8'd 591  ;
mem[ 592 ]=8'd 592  ;
mem[ 593 ]=8'd 593  ;
mem[ 594 ]=8'd 594  ;
mem[ 595 ]=8'd 595  ;
mem[ 596 ]=8'd 596  ;
mem[ 597 ]=8'd 597  ;
mem[ 598 ]=8'd 598  ;
mem[ 599 ]=8'd 599  ;
mem[ 600 ]=8'd 600  ;
mem[ 601 ]=8'd 601  ;
mem[ 602 ]=8'd 602  ;
mem[ 603 ]=8'd 603  ;
mem[ 604 ]=8'd 604  ;
mem[ 605 ]=8'd 605  ;
mem[ 606 ]=8'd 606  ;
mem[ 607 ]=8'd 607  ;
mem[ 608 ]=8'd 608  ;
mem[ 609 ]=8'd 609  ;
mem[ 610 ]=8'd 610  ;
mem[ 611 ]=8'd 611  ;
mem[ 612 ]=8'd 612  ;
mem[ 613 ]=8'd 613  ;
mem[ 614 ]=8'd 614  ;
mem[ 615 ]=8'd 615  ;
mem[ 616 ]=8'd 616  ;
mem[ 617 ]=8'd 617  ;
mem[ 618 ]=8'd 618  ;
mem[ 619 ]=8'd 619  ;
mem[ 620 ]=8'd 620  ;
mem[ 621 ]=8'd 621  ;
mem[ 622 ]=8'd 622  ;
mem[ 623 ]=8'd 623  ;
mem[ 624 ]=8'd 624  ;
mem[ 625 ]=8'd 625  ;
mem[ 626 ]=8'd 626  ;
mem[ 627 ]=8'd 627  ;
mem[ 628 ]=8'd 628  ;
mem[ 629 ]=8'd 629  ;
mem[ 630 ]=8'd 630  ;
mem[ 631 ]=8'd 631  ;
mem[ 632 ]=8'd 632  ;
mem[ 633 ]=8'd 633  ;
mem[ 634 ]=8'd 634  ;
mem[ 635 ]=8'd 635  ;
mem[ 636 ]=8'd 636  ;
mem[ 637 ]=8'd 637  ;
mem[ 638 ]=8'd 638  ;
mem[ 639 ]=8'd 639  ;
mem[ 640 ]=8'd 640  ;
mem[ 641 ]=8'd 641  ;
mem[ 642 ]=8'd 642  ;
mem[ 643 ]=8'd 643  ;
mem[ 644 ]=8'd 644  ;
mem[ 645 ]=8'd 645  ;
mem[ 646 ]=8'd 646  ;
mem[ 647 ]=8'd 647  ;
mem[ 648 ]=8'd 648  ;
mem[ 649 ]=8'd 649  ;
mem[ 650 ]=8'd 650  ;
mem[ 651 ]=8'd 651  ;
mem[ 652 ]=8'd 652  ;
mem[ 653 ]=8'd 653  ;
mem[ 654 ]=8'd 654  ;
mem[ 655 ]=8'd 655  ;
mem[ 656 ]=8'd 656  ;
mem[ 657 ]=8'd 657  ;
mem[ 658 ]=8'd 658  ;
mem[ 659 ]=8'd 659  ;
mem[ 660 ]=8'd 660  ;
mem[ 661 ]=8'd 661  ;
mem[ 662 ]=8'd 662  ;
mem[ 663 ]=8'd 663  ;
mem[ 664 ]=8'd 664  ;
mem[ 665 ]=8'd 665  ;
mem[ 666 ]=8'd 666  ;
mem[ 667 ]=8'd 667  ;
mem[ 668 ]=8'd 668  ;
mem[ 669 ]=8'd 669  ;
mem[ 670 ]=8'd 670  ;
mem[ 671 ]=8'd 671  ;
mem[ 672 ]=8'd 672  ;
mem[ 673 ]=8'd 673  ;
mem[ 674 ]=8'd 674  ;
mem[ 675 ]=8'd 675  ;
mem[ 676 ]=8'd 676  ;
mem[ 677 ]=8'd 677  ;
mem[ 678 ]=8'd 678  ;
mem[ 679 ]=8'd 679  ;
mem[ 680 ]=8'd 680  ;
mem[ 681 ]=8'd 681  ;
mem[ 682 ]=8'd 682  ;
mem[ 683 ]=8'd 683  ;
mem[ 684 ]=8'd 684  ;
mem[ 685 ]=8'd 685  ;
mem[ 686 ]=8'd 686  ;
mem[ 687 ]=8'd 687  ;
mem[ 688 ]=8'd 688  ;
mem[ 689 ]=8'd 689  ;
mem[ 690 ]=8'd 690  ;
mem[ 691 ]=8'd 691  ;
mem[ 692 ]=8'd 692  ;
mem[ 693 ]=8'd 693  ;
mem[ 694 ]=8'd 694  ;
mem[ 695 ]=8'd 695  ;
mem[ 696 ]=8'd 696  ;
mem[ 697 ]=8'd 697  ;
mem[ 698 ]=8'd 698  ;
mem[ 699 ]=8'd 699  ;
mem[ 700 ]=8'd 700  ;
mem[ 701 ]=8'd 701  ;
mem[ 702 ]=8'd 702  ;
mem[ 703 ]=8'd 703  ;
mem[ 704 ]=8'd 704  ;
mem[ 705 ]=8'd 705  ;
mem[ 706 ]=8'd 706  ;
mem[ 707 ]=8'd 707  ;
mem[ 708 ]=8'd 708  ;
mem[ 709 ]=8'd 709  ;
mem[ 710 ]=8'd 710  ;
mem[ 711 ]=8'd 711  ;
mem[ 712 ]=8'd 712  ;
mem[ 713 ]=8'd 713  ;
mem[ 714 ]=8'd 714  ;
mem[ 715 ]=8'd 715  ;
mem[ 716 ]=8'd 716  ;
mem[ 717 ]=8'd 717  ;
mem[ 718 ]=8'd 718  ;
mem[ 719 ]=8'd 719  ;
mem[ 720 ]=8'd 720  ;
mem[ 721 ]=8'd 721  ;
mem[ 722 ]=8'd 722  ;
mem[ 723 ]=8'd 723  ;
mem[ 724 ]=8'd 724  ;
mem[ 725 ]=8'd 725  ;
mem[ 726 ]=8'd 726  ;
mem[ 727 ]=8'd 727  ;
mem[ 728 ]=8'd 728  ;
mem[ 729 ]=8'd 729  ;
mem[ 730 ]=8'd 730  ;
mem[ 731 ]=8'd 731  ;
mem[ 732 ]=8'd 732  ;
mem[ 733 ]=8'd 733  ;
mem[ 734 ]=8'd 734  ;
mem[ 735 ]=8'd 735  ;
mem[ 736 ]=8'd 736  ;
mem[ 737 ]=8'd 737  ;
mem[ 738 ]=8'd 738  ;
mem[ 739 ]=8'd 739  ;
mem[ 740 ]=8'd 740  ;
mem[ 741 ]=8'd 741  ;
mem[ 742 ]=8'd 742  ;
mem[ 743 ]=8'd 743  ;
mem[ 744 ]=8'd 744  ;
mem[ 745 ]=8'd 745  ;
mem[ 746 ]=8'd 746  ;
mem[ 747 ]=8'd 747  ;
mem[ 748 ]=8'd 748  ;
mem[ 749 ]=8'd 749  ;
mem[ 750 ]=8'd 750  ;
mem[ 751 ]=8'd 751  ;
mem[ 752 ]=8'd 752  ;
mem[ 753 ]=8'd 753  ;
mem[ 754 ]=8'd 754  ;
mem[ 755 ]=8'd 755  ;
mem[ 756 ]=8'd 756  ;
mem[ 757 ]=8'd 757  ;
mem[ 758 ]=8'd 758  ;
mem[ 759 ]=8'd 759  ;
mem[ 760 ]=8'd 760  ;
mem[ 761 ]=8'd 761  ;
mem[ 762 ]=8'd 762  ;
mem[ 763 ]=8'd 763  ;
mem[ 764 ]=8'd 764  ;
mem[ 765 ]=8'd 765  ;
mem[ 766 ]=8'd 766  ;
mem[ 767 ]=8'd 767  ;
mem[ 768 ]=8'd 768  ;
mem[ 769 ]=8'd 769  ;
mem[ 770 ]=8'd 770  ;
mem[ 771 ]=8'd 771  ;
mem[ 772 ]=8'd 772  ;
mem[ 773 ]=8'd 773  ;
mem[ 774 ]=8'd 774  ;
mem[ 775 ]=8'd 775  ;
mem[ 776 ]=8'd 776  ;
mem[ 777 ]=8'd 777  ;
mem[ 778 ]=8'd 778  ;
mem[ 779 ]=8'd 779  ;
mem[ 780 ]=8'd 780  ;
mem[ 781 ]=8'd 781  ;
mem[ 782 ]=8'd 782  ;
mem[ 783 ]=8'd 783  ;
mem[ 784 ]=8'd 784  ;
mem[ 785 ]=8'd 785  ;
mem[ 786 ]=8'd 786  ;
mem[ 787 ]=8'd 787  ;
mem[ 788 ]=8'd 788  ;
mem[ 789 ]=8'd 789  ;
mem[ 790 ]=8'd 790  ;
mem[ 791 ]=8'd 791  ;
mem[ 792 ]=8'd 792  ;
mem[ 793 ]=8'd 793  ;
mem[ 794 ]=8'd 794  ;
mem[ 795 ]=8'd 795  ;
mem[ 796 ]=8'd 796  ;
mem[ 797 ]=8'd 797  ;
mem[ 798 ]=8'd 798  ;
mem[ 799 ]=8'd 799  ;
mem[ 800 ]=8'd 800  ;
mem[ 801 ]=8'd 801  ;
mem[ 802 ]=8'd 802  ;
mem[ 803 ]=8'd 803  ;
mem[ 804 ]=8'd 804  ;
mem[ 805 ]=8'd 805  ;
mem[ 806 ]=8'd 806  ;
mem[ 807 ]=8'd 807  ;
mem[ 808 ]=8'd 808  ;
mem[ 809 ]=8'd 809  ;
mem[ 810 ]=8'd 810  ;
mem[ 811 ]=8'd 811  ;
mem[ 812 ]=8'd 812  ;
mem[ 813 ]=8'd 813  ;
mem[ 814 ]=8'd 814  ;
mem[ 815 ]=8'd 815  ;
mem[ 816 ]=8'd 816  ;
mem[ 817 ]=8'd 817  ;
mem[ 818 ]=8'd 818  ;
mem[ 819 ]=8'd 819  ;
mem[ 820 ]=8'd 820  ;
mem[ 821 ]=8'd 821  ;
mem[ 822 ]=8'd 822  ;
mem[ 823 ]=8'd 823  ;
mem[ 824 ]=8'd 824  ;
mem[ 825 ]=8'd 825  ;
mem[ 826 ]=8'd 826  ;
mem[ 827 ]=8'd 827  ;
mem[ 828 ]=8'd 828  ;
mem[ 829 ]=8'd 829  ;
mem[ 830 ]=8'd 830  ;
mem[ 831 ]=8'd 831  ;
mem[ 832 ]=8'd 832  ;
mem[ 833 ]=8'd 833  ;
mem[ 834 ]=8'd 834  ;
mem[ 835 ]=8'd 835  ;
mem[ 836 ]=8'd 836  ;
mem[ 837 ]=8'd 837  ;
mem[ 838 ]=8'd 838  ;
mem[ 839 ]=8'd 839  ;
mem[ 840 ]=8'd 840  ;
mem[ 841 ]=8'd 841  ;
mem[ 842 ]=8'd 842  ;
mem[ 843 ]=8'd 843  ;
mem[ 844 ]=8'd 844  ;
mem[ 845 ]=8'd 845  ;
mem[ 846 ]=8'd 846  ;
mem[ 847 ]=8'd 847  ;
mem[ 848 ]=8'd 848  ;
mem[ 849 ]=8'd 849  ;
mem[ 850 ]=8'd 850  ;
mem[ 851 ]=8'd 851  ;
mem[ 852 ]=8'd 852  ;
mem[ 853 ]=8'd 853  ;
mem[ 854 ]=8'd 854  ;
mem[ 855 ]=8'd 855  ;
mem[ 856 ]=8'd 856  ;
mem[ 857 ]=8'd 857  ;
mem[ 858 ]=8'd 858  ;
mem[ 859 ]=8'd 859  ;
mem[ 860 ]=8'd 860  ;
mem[ 861 ]=8'd 861  ;
mem[ 862 ]=8'd 862  ;
mem[ 863 ]=8'd 863  ;
mem[ 864 ]=8'd 864  ;
mem[ 865 ]=8'd 865  ;
mem[ 866 ]=8'd 866  ;
mem[ 867 ]=8'd 867  ;
mem[ 868 ]=8'd 868  ;
mem[ 869 ]=8'd 869  ;
mem[ 870 ]=8'd 870  ;
mem[ 871 ]=8'd 871  ;
mem[ 872 ]=8'd 872  ;
mem[ 873 ]=8'd 873  ;
mem[ 874 ]=8'd 874  ;
mem[ 875 ]=8'd 875  ;
mem[ 876 ]=8'd 876  ;
mem[ 877 ]=8'd 877  ;
mem[ 878 ]=8'd 878  ;
mem[ 879 ]=8'd 879  ;
mem[ 880 ]=8'd 880  ;
mem[ 881 ]=8'd 881  ;
mem[ 882 ]=8'd 882  ;
mem[ 883 ]=8'd 883  ;
mem[ 884 ]=8'd 884  ;
mem[ 885 ]=8'd 885  ;
mem[ 886 ]=8'd 886  ;
mem[ 887 ]=8'd 887  ;
mem[ 888 ]=8'd 888  ;
mem[ 889 ]=8'd 889  ;
mem[ 890 ]=8'd 890  ;
mem[ 891 ]=8'd 891  ;
mem[ 892 ]=8'd 892  ;
mem[ 893 ]=8'd 893  ;
mem[ 894 ]=8'd 894  ;
mem[ 895 ]=8'd 895  ;
mem[ 896 ]=8'd 896  ;
mem[ 897 ]=8'd 897  ;
mem[ 898 ]=8'd 898  ;
mem[ 899 ]=8'd 899  ;
mem[ 900 ]=8'd 900  ;
mem[ 901 ]=8'd 901  ;
mem[ 902 ]=8'd 902  ;
mem[ 903 ]=8'd 903  ;
mem[ 904 ]=8'd 904  ;
mem[ 905 ]=8'd 905  ;
mem[ 906 ]=8'd 906  ;
mem[ 907 ]=8'd 907  ;
mem[ 908 ]=8'd 908  ;
mem[ 909 ]=8'd 909  ;
mem[ 910 ]=8'd 910  ;
mem[ 911 ]=8'd 911  ;
mem[ 912 ]=8'd 912  ;
mem[ 913 ]=8'd 913  ;
mem[ 914 ]=8'd 914  ;
mem[ 915 ]=8'd 915  ;
mem[ 916 ]=8'd 916  ;
mem[ 917 ]=8'd 917  ;
mem[ 918 ]=8'd 918  ;
mem[ 919 ]=8'd 919  ;
mem[ 920 ]=8'd 920  ;
mem[ 921 ]=8'd 921  ;
mem[ 922 ]=8'd 922  ;
mem[ 923 ]=8'd 923  ;
mem[ 924 ]=8'd 924  ;
mem[ 925 ]=8'd 925  ;
mem[ 926 ]=8'd 926  ;
mem[ 927 ]=8'd 927  ;
mem[ 928 ]=8'd 928  ;
mem[ 929 ]=8'd 929  ;
mem[ 930 ]=8'd 930  ;
mem[ 931 ]=8'd 931  ;
mem[ 932 ]=8'd 932  ;
mem[ 933 ]=8'd 933  ;
mem[ 934 ]=8'd 934  ;
mem[ 935 ]=8'd 935  ;
mem[ 936 ]=8'd 936  ;
mem[ 937 ]=8'd 937  ;
mem[ 938 ]=8'd 938  ;
mem[ 939 ]=8'd 939  ;
mem[ 940 ]=8'd 940  ;
mem[ 941 ]=8'd 941  ;
mem[ 942 ]=8'd 942  ;
mem[ 943 ]=8'd 943  ;
mem[ 944 ]=8'd 944  ;
mem[ 945 ]=8'd 945  ;
mem[ 946 ]=8'd 946  ;
mem[ 947 ]=8'd 947  ;
mem[ 948 ]=8'd 948  ;
mem[ 949 ]=8'd 949  ;
mem[ 950 ]=8'd 950  ;
mem[ 951 ]=8'd 951  ;
mem[ 952 ]=8'd 952  ;
mem[ 953 ]=8'd 953  ;
mem[ 954 ]=8'd 954  ;
mem[ 955 ]=8'd 955  ;
mem[ 956 ]=8'd 956  ;
mem[ 957 ]=8'd 957  ;
mem[ 958 ]=8'd 958  ;
mem[ 959 ]=8'd 959  ;
mem[ 960 ]=8'd 960  ;
mem[ 961 ]=8'd 961  ;
mem[ 962 ]=8'd 962  ;
mem[ 963 ]=8'd 963  ;
mem[ 964 ]=8'd 964  ;
mem[ 965 ]=8'd 965  ;
mem[ 966 ]=8'd 966  ;
mem[ 967 ]=8'd 967  ;
mem[ 968 ]=8'd 968  ;
mem[ 969 ]=8'd 969  ;
mem[ 970 ]=8'd 970  ;
mem[ 971 ]=8'd 971  ;
mem[ 972 ]=8'd 972  ;
mem[ 973 ]=8'd 973  ;
mem[ 974 ]=8'd 974  ;
mem[ 975 ]=8'd 975  ;
mem[ 976 ]=8'd 976  ;
mem[ 977 ]=8'd 977  ;
mem[ 978 ]=8'd 978  ;
mem[ 979 ]=8'd 979  ;
mem[ 980 ]=8'd 980  ;
mem[ 981 ]=8'd 981  ;
mem[ 982 ]=8'd 982  ;
mem[ 983 ]=8'd 983  ;
mem[ 984 ]=8'd 984  ;
mem[ 985 ]=8'd 985  ;
mem[ 986 ]=8'd 986  ;
mem[ 987 ]=8'd 987  ;
mem[ 988 ]=8'd 988  ;
mem[ 989 ]=8'd 989  ;
mem[ 990 ]=8'd 990  ;
mem[ 991 ]=8'd 991  ;
mem[ 992 ]=8'd 992  ;
mem[ 993 ]=8'd 993  ;
mem[ 994 ]=8'd 994  ;
mem[ 995 ]=8'd 995  ;
mem[ 996 ]=8'd 996  ;
mem[ 997 ]=8'd 997  ;
mem[ 998 ]=8'd 998  ;
mem[ 999 ]=8'd 999  ;
mem[ 1000 ]=8'd 1000  ;
mem[ 1001 ]=8'd 1001  ;
mem[ 1002 ]=8'd 1002  ;
mem[ 1003 ]=8'd 1003  ;
mem[ 1004 ]=8'd 1004  ;
mem[ 1005 ]=8'd 1005  ;
mem[ 1006 ]=8'd 1006  ;
mem[ 1007 ]=8'd 1007  ;
mem[ 1008 ]=8'd 1008  ;
mem[ 1009 ]=8'd 1009  ;
mem[ 1010 ]=8'd 1010  ;
mem[ 1011 ]=8'd 1011  ;
mem[ 1012 ]=8'd 1012  ;
mem[ 1013 ]=8'd 1013  ;
mem[ 1014 ]=8'd 1014  ;
mem[ 1015 ]=8'd 1015  ;
mem[ 1016 ]=8'd 1016  ;
mem[ 1017 ]=8'd 1017  ;
mem[ 1018 ]=8'd 1018  ;
mem[ 1019 ]=8'd 1019  ;
mem[ 1020 ]=8'd 1020  ;
mem[ 1021 ]=8'd 1021  ;
mem[ 1022 ]=8'd 1022  ;
mem[ 1023 ]=8'd 1023  ;
end

            
        
	 
	 
	 
	 
endmodule
